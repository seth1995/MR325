#test
R1 0 1  1
C1 1 2  1
C2 1 0  1
Vin 2 0  0 sin 1 2 2500M 0
.tran TR 0 1n 1p
.end