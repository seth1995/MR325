#a circuit has diode
MP1 2 1 3 4 1
MN1 2 1 0 2 1
V1 1 0 1.7
V2 3 0 1.7

.end