*NOR
MP1 4 1 5 4 1
MP2 3 2 4 4 1
MN1 3 2 0 2 1
MN2 3 1 0 2 1
VDD 5 0 3
VA 1 0 0 pulse 0.7 2.2 1n 1n 20n 30n
VB 2 0 0 pulse 0.7 2.2 1n 1n 20n 30n
C1 3 0 0.003p
.tran TR 0 100n 100p
.END