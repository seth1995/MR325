* mosfet off A w o-
Vin 1 0 0.7 
Vdd 2 0 1.8
C1 2 0 1p
MP1 3 1 2 4 1
MN1 3 1 0 2 1

.TRAN TR 0 10u 5u
.END
