*NAND
MP1 4 1 3 4 1
MP2 4 2 3 4 1
MN1 4 1 5 2 1
MN2 5 2 0 2 1
VDD 3 0 3
VA 1 0 0 pulse 0 3 1n 1n 20n 30n
VB 2 0 0 pulse 3 0 1n 1n 20n 30n
C1 4 0 0.003p
.tran TR 0 100n 100p
.END