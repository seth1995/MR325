*acMOS

V1 1 0 5 
R1 1 2 5

C3 2 0 0.2
L1 1 2 0.1


.AC DEC 10 0.01 10k
.END