*ac CL
V1 1 0 1
R1 1 2 5MEG
C1 2 0 0.2u
.AC DEC 10 0.01 10

.END