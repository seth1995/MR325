* buffer
* Vin 1 0 0 sin 1.5 1.5 80M 0
Vin 1 0 1	pulse 3 0 0 0 20n 30n
Vdd 2 0 3
C1 3 0 1p
MP2 3 1 2 40 1
MN1 3 1 0 20 1

C2 5 0 10p
MP3 5 3 2 40 1
MN4 5 3 0 20 1



C3 7 0 10p
MP5 7 5 2 40 1
MN6 7 5 0 20 1



C4 8 0 10p
MP7 8 7 2 40 1
MN8 8 7 0 20 1



C5 9 0 10p
MP9  9 8 2 40 1
MN10  9 8 0 20 1

C6 10 0 10p
MP11 10 9 2 40 1
MN12 10 9 0 20 1



C7 11 0 10p
MP13  11 10 2 40 1
MN14  11 10 0 20 1

C8 12 0 10p
MP15 12 11 2 40 1
MN16 12 11 0 20 1




C9 13 0 10p
MP13  13 12 2 40 1
MN14  13 12 0 20 1

C10 14 0 10p
MP15 14 13 2 40 1
MN16 14 13 0 20 1



C11 15 0 10p
MP13  15 14 2 40 1
MN14  15 14 0 20 1

C12 16 0 10p
MP15 16 15 2 40 1
MN16 16 15 0 20 1

*.DC  Vin 0 3 0.01
.tran TR 0 100n 10p
.END

