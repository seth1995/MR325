* tran1
V1 1 0 5
R2 1 2 5
C3 2 0 0.2

.TRAN TR 0 10 0.001
.END